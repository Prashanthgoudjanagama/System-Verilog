
// file name : 18_practive_fork_join.sv
// module name : top_practive_fork_join

